library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use IEEE.NUMERIC_STD.ALL;

entity conv_layer_1 is
    Port (
        w : in STD_LOGIC_VECTOR (3*3*3-1 downto 0);
        x : in STD_LOGIC_VECTOR (32*32*3*8-1 downto 0);
        cnt : in STD_LOGIC_VECTOR(9 downto 0);
        --done : out STD_LOGIC;
        z : out STD_LOGIC_VECTOR (14 downto 0)
        );
end conv_layer_1;

architecture Behavioral of conv_layer_1 is
    component single_step_conv_1
            Port ( 
                    w : in STD_LOGIC_VECTOR (3*3*3-1 downto 0);
                    x : in STD_LOGIC_VECTOR (3*3*3*8-1 downto 0);
                    c : in STD_LOGIC_VECTOR (3 downto 0);
                    z : out STD_LOGIC_VECTOR (14 downto 0)
                 );
    end component;

    
    signal S : STD_LOGIC_VECTOR(9 downto 0) := (others => '0');--conv state 
    signal x_single : STD_LOGIC_VECTOR(3*3*3*8-1 downto 0);--input for single step conv
    signal c : STD_LOGIC_VECTOR (3 downto 0);
    signal z_single : STD_LOGIC_VECTOR(14 downto 0);
begin

    z <= z_single;                      

    uut: single_step_conv_1 port map ( --w => weight,
                                     w => w,
                                     x => x_single,
                                     c => c,
                                     z => z_single
                                    );

    --S <= cnt(9 downto 6) & cnt(1) & cnt(5 downto 2) & cnt(0);--order of output for next pooling layer
    S <= cnt(9 downto 0);
    
    L1: for m in 0 to 2 generate 
        process(S, x)
            variable I : integer;
        begin
            I := to_integer(unsigned(S));
            case(S) is
                when "0000000000" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= x(32*32*m*8+33*8+7 downto 32*32*m*8+32*8) & "00000000" & x(32*32*m*8+1*8+7 downto 32*32*m*8) & "00000000000000000000000000000000";--p0 the left top corner

                when "0000000001" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= x(32*32*m*8+34*8+7 downto 32*32*m*8+32*8) & x(32*32*m*8+2*8+7 downto 32*32*m*8) & "000000000000000000000000";--p1 the top edge
                when "0000000010" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= x(32*32*m*8+35*8+7 downto 32*32*m*8+33*8) & x(32*32*m*8+3*8+7 downto 32*32*m*8+1*8) & "000000000000000000000000";
                when "0000000011" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= x(32*32*m*8+36*8+7 downto 32*32*m*8+34*8) & x(32*32*m*8+4*8+7 downto 32*32*m*8+2*8) & "000000000000000000000000";
                when "0000000100" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= x(32*32*m*8+37*8+7 downto 32*32*m*8+35*8) & x(32*32*m*8+5*8+7 downto 32*32*m*8+3*8) & "000000000000000000000000";
                when "0000000101" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= x(32*32*m*8+38*8+7 downto 32*32*m*8+36*8) & x(32*32*m*8+6*8+7 downto 32*32*m*8+4*8) & "000000000000000000000000";
                when "0000000110" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= x(32*32*m*8+39*8+7 downto 32*32*m*8+37*8) & x(32*32*m*8+7*8+7 downto 32*32*m*8+5*8) & "000000000000000000000000";
                when "0000000111" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= x(32*32*m*8+40*8+7 downto 32*32*m*8+38*8) & x(32*32*m*8+8*8+7 downto 32*32*m*8+6*8) & "000000000000000000000000";
                when "0000001000" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= x(32*32*m*8+41*8+7 downto 32*32*m*8+39*8) & x(32*32*m*8+9*8+7 downto 32*32*m*8+7*8) & "000000000000000000000000";
                when "0000001001" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= x(32*32*m*8+42*8+7 downto 32*32*m*8+40*8) & x(32*32*m*8+10*8+7 downto 32*32*m*8+8*8) & "000000000000000000000000";
                when "0000001010" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= x(32*32*m*8+43*8+7 downto 32*32*m*8+41*8) & x(32*32*m*8+11*8+7 downto 32*32*m*8+9*8) & "000000000000000000000000";
                when "0000001011" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= x(32*32*m*8+44*8+7 downto 32*32*m*8+42*8) & x(32*32*m*8+12*8+7 downto 32*32*m*8+10*8) & "000000000000000000000000";
                when "0000001100" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= x(32*32*m*8+45*8+7 downto 32*32*m*8+43*8) & x(32*32*m*8+13*8+7 downto 32*32*m*8+11*8) & "000000000000000000000000";
                when "0000001101" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= x(32*32*m*8+46*8+7 downto 32*32*m*8+44*8) & x(32*32*m*8+14*8+7 downto 32*32*m*8+12*8) & "000000000000000000000000";
                when "0000001110" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= x(32*32*m*8+47*8+7 downto 32*32*m*8+45*8) & x(32*32*m*8+15*8+7 downto 32*32*m*8+13*8) & "000000000000000000000000";
                when "0000001111" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= x(32*32*m*8+48*8+7 downto 32*32*m*8+46*8) & x(32*32*m*8+16*8+7 downto 32*32*m*8+14*8) & "000000000000000000000000";
                when "0000010000" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= x(32*32*m*8+49*8+7 downto 32*32*m*8+47*8) & x(32*32*m*8+17*8+7 downto 32*32*m*8+15*8) & "000000000000000000000000";
                when "0000010001" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= x(32*32*m*8+50*8+7 downto 32*32*m*8+48*8) & x(32*32*m*8+18*8+7 downto 32*32*m*8+16*8) & "000000000000000000000000";
                when "0000010010" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= x(32*32*m*8+51*8+7 downto 32*32*m*8+49*8) & x(32*32*m*8+19*8+7 downto 32*32*m*8+17*8) & "000000000000000000000000";
                when "0000010011" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= x(32*32*m*8+52*8+7 downto 32*32*m*8+50*8) & x(32*32*m*8+20*8+7 downto 32*32*m*8+18*8) & "000000000000000000000000";
                when "0000010100" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= x(32*32*m*8+53*8+7 downto 32*32*m*8+51*8) & x(32*32*m*8+21*8+7 downto 32*32*m*8+19*8) & "000000000000000000000000";
                when "0000010101" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= x(32*32*m*8+54*8+7 downto 32*32*m*8+52*8) & x(32*32*m*8+22*8+7 downto 32*32*m*8+20*8) & "000000000000000000000000";
                when "0000010110" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= x(32*32*m*8+55*8+7 downto 32*32*m*8+53*8) & x(32*32*m*8+23*8+7 downto 32*32*m*8+21*8) & "000000000000000000000000";
                when "0000010111" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= x(32*32*m*8+56*8+7 downto 32*32*m*8+54*8) & x(32*32*m*8+24*8+7 downto 32*32*m*8+22*8) & "000000000000000000000000";
                when "0000011000" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= x(32*32*m*8+57*8+7 downto 32*32*m*8+55*8) & x(32*32*m*8+25*8+7 downto 32*32*m*8+23*8) & "000000000000000000000000";
                when "0000011001" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= x(32*32*m*8+58*8+7 downto 32*32*m*8+56*8) & x(32*32*m*8+26*8+7 downto 32*32*m*8+24*8) & "000000000000000000000000";
                when "0000011010" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= x(32*32*m*8+59*8+7 downto 32*32*m*8+57*8) & x(32*32*m*8+27*8+7 downto 32*32*m*8+25*8) & "000000000000000000000000";
                when "0000011011" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= x(32*32*m*8+60*8+7 downto 32*32*m*8+58*8) & x(32*32*m*8+28*8+7 downto 32*32*m*8+26*8) & "000000000000000000000000";
                when "0000011100" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= x(32*32*m*8+61*8+7 downto 32*32*m*8+59*8) & x(32*32*m*8+29*8+7 downto 32*32*m*8+27*8) & "000000000000000000000000";
                when "0000011101" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= x(32*32*m*8+62*8+7 downto 32*32*m*8+60*8) & x(32*32*m*8+30*8+7 downto 32*32*m*8+28*8) & "000000000000000000000000";
                when "0000011110" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= x(32*32*m*8+63*8+7 downto 32*32*m*8+61*8) & x(32*32*m*8+31*8+7 downto 32*32*m*8+29*8) & "000000000000000000000000";

                when "0000011111" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= "00000000" & x(32*32*m*8+63*8+7 downto 32*32*m*8+62*8) & "00000000" & x(32*32*m*8+31*8+7 downto 32*32*m*8+30*8) & "000000000000000000000000";--p2 the right top corner

                when "0000100000" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= x(32*32*m*8+65*8+7 downto 32*32*m*8+64*8) & "00000000" & x(32*32*m*8+33*8+7 downto 32*32*m*8+32*8) & "00000000" & x(32*32*m*8+1*8+7 downto 32*32*m*8) & "00000000";--p3 the left edge
                when "0001000000" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= x(32*32*m*8+97*8+7 downto 32*32*m*8+96*8) & "00000000" & x(32*32*m*8+65*8+7 downto 32*32*m*8+64*8) & "00000000" & x(32*32*m*8+33*8+7 downto 32*32*m*8+32*8) & "00000000";
                when "0001100000" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= x(32*32*m*8+129*8+7 downto 32*32*m*8+128*8) & "00000000" & x(32*32*m*8+97*8+7 downto 32*32*m*8+96*8) & "00000000" & x(32*32*m*8+65*8+7 downto 32*32*m*8+64*8) & "00000000";
                when "0010000000" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= x(32*32*m*8+161*8+7 downto 32*32*m*8+160*8) & "00000000" & x(32*32*m*8+129*8+7 downto 32*32*m*8+128*8) & "00000000" & x(32*32*m*8+97*8+7 downto 32*32*m*8+96*8) & "00000000";
                when "0010100000" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= x(32*32*m*8+193*8+7 downto 32*32*m*8+192*8) & "00000000" & x(32*32*m*8+161*8+7 downto 32*32*m*8+160*8) & "00000000" & x(32*32*m*8+129*8+7 downto 32*32*m*8+128*8) & "00000000";
                when "0011000000" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= x(32*32*m*8+225*8+7 downto 32*32*m*8+224*8) & "00000000" & x(32*32*m*8+193*8+7 downto 32*32*m*8+192*8) & "00000000" & x(32*32*m*8+161*8+7 downto 32*32*m*8+160*8) & "00000000";
                when "0011100000" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= x(32*32*m*8+257*8+7 downto 32*32*m*8+256*8) & "00000000" & x(32*32*m*8+225*8+7 downto 32*32*m*8+224*8) & "00000000" & x(32*32*m*8+193*8+7 downto 32*32*m*8+192*8) & "00000000";
                when "0100000000" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= x(32*32*m*8+289*8+7 downto 32*32*m*8+288*8) & "00000000" & x(32*32*m*8+257*8+7 downto 32*32*m*8+256*8) & "00000000" & x(32*32*m*8+225*8+7 downto 32*32*m*8+224*8) & "00000000";
                when "0100100000" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= x(32*32*m*8+321*8+7 downto 32*32*m*8+320*8) & "00000000" & x(32*32*m*8+289*8+7 downto 32*32*m*8+288*8) & "00000000" & x(32*32*m*8+257*8+7 downto 32*32*m*8+256*8) & "00000000";
                when "0101000000" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= x(32*32*m*8+353*8+7 downto 32*32*m*8+352*8) & "00000000" & x(32*32*m*8+321*8+7 downto 32*32*m*8+320*8) & "00000000" & x(32*32*m*8+289*8+7 downto 32*32*m*8+288*8) & "00000000";
                when "0101100000" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= x(32*32*m*8+385*8+7 downto 32*32*m*8+384*8) & "00000000" & x(32*32*m*8+353*8+7 downto 32*32*m*8+352*8) & "00000000" & x(32*32*m*8+321*8+7 downto 32*32*m*8+320*8) & "00000000";
                when "0110000000" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= x(32*32*m*8+417*8+7 downto 32*32*m*8+416*8) & "00000000" & x(32*32*m*8+385*8+7 downto 32*32*m*8+384*8) & "00000000" & x(32*32*m*8+353*8+7 downto 32*32*m*8+352*8) & "00000000";
                when "0110100000" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= x(32*32*m*8+449*8+7 downto 32*32*m*8+448*8) & "00000000" & x(32*32*m*8+417*8+7 downto 32*32*m*8+416*8) & "00000000" & x(32*32*m*8+385*8+7 downto 32*32*m*8+384*8) & "00000000";
                when "0111000000" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= x(32*32*m*8+481*8+7 downto 32*32*m*8+480*8) & "00000000" & x(32*32*m*8+449*8+7 downto 32*32*m*8+448*8) & "00000000" & x(32*32*m*8+417*8+7 downto 32*32*m*8+416*8) & "00000000";
                when "0111100000" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= x(32*32*m*8+513*8+7 downto 32*32*m*8+512*8) & "00000000" & x(32*32*m*8+481*8+7 downto 32*32*m*8+480*8) & "00000000" & x(32*32*m*8+449*8+7 downto 32*32*m*8+448*8) & "00000000";
                when "1000000000" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= x(32*32*m*8+545*8+7 downto 32*32*m*8+544*8) & "00000000" & x(32*32*m*8+513*8+7 downto 32*32*m*8+512*8) & "00000000" & x(32*32*m*8+481*8+7 downto 32*32*m*8+480*8) & "00000000";
                when "1000100000" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= x(32*32*m*8+577*8+7 downto 32*32*m*8+576*8) & "00000000" & x(32*32*m*8+545*8+7 downto 32*32*m*8+544*8) & "00000000" & x(32*32*m*8+513*8+7 downto 32*32*m*8+512*8) & "00000000";
                when "1001000000" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= x(32*32*m*8+609*8+7 downto 32*32*m*8+608*8) & "00000000" & x(32*32*m*8+577*8+7 downto 32*32*m*8+576*8) & "00000000" & x(32*32*m*8+545*8+7 downto 32*32*m*8+544*8) & "00000000";
                when "1001100000" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= x(32*32*m*8+641*8+7 downto 32*32*m*8+640*8) & "00000000" & x(32*32*m*8+609*8+7 downto 32*32*m*8+608*8) & "00000000" & x(32*32*m*8+577*8+7 downto 32*32*m*8+576*8) & "00000000";
                when "1010000000" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= x(32*32*m*8+673*8+7 downto 32*32*m*8+672*8) & "00000000" & x(32*32*m*8+641*8+7 downto 32*32*m*8+640*8) & "00000000" & x(32*32*m*8+609*8+7 downto 32*32*m*8+608*8) & "00000000";
                when "1010100000" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= x(32*32*m*8+705*8+7 downto 32*32*m*8+704*8) & "00000000" & x(32*32*m*8+673*8+7 downto 32*32*m*8+672*8) & "00000000" & x(32*32*m*8+641*8+7 downto 32*32*m*8+640*8) & "00000000";
                when "1011000000" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= x(32*32*m*8+737*8+7 downto 32*32*m*8+736*8) & "00000000" & x(32*32*m*8+705*8+7 downto 32*32*m*8+704*8) & "00000000" & x(32*32*m*8+673*8+7 downto 32*32*m*8+672*8) & "00000000";
                when "1011100000" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= x(32*32*m*8+769*8+7 downto 32*32*m*8+768*8) & "00000000" & x(32*32*m*8+737*8+7 downto 32*32*m*8+736*8) & "00000000" & x(32*32*m*8+705*8+7 downto 32*32*m*8+704*8) & "00000000";
                when "1100000000" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= x(32*32*m*8+801*8+7 downto 32*32*m*8+800*8) & "00000000" & x(32*32*m*8+769*8+7 downto 32*32*m*8+768*8) & "00000000" & x(32*32*m*8+737*8+7 downto 32*32*m*8+736*8) & "00000000";
                when "1100100000" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= x(32*32*m*8+833*8+7 downto 32*32*m*8+832*8) & "00000000" & x(32*32*m*8+801*8+7 downto 32*32*m*8+800*8) & "00000000" & x(32*32*m*8+769*8+7 downto 32*32*m*8+768*8) & "00000000";
                when "1101000000" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= x(32*32*m*8+865*8+7 downto 32*32*m*8+864*8) & "00000000" & x(32*32*m*8+833*8+7 downto 32*32*m*8+832*8) & "00000000" & x(32*32*m*8+801*8+7 downto 32*32*m*8+800*8) & "00000000";
                when "1101100000" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= x(32*32*m*8+897*8+7 downto 32*32*m*8+896*8) & "00000000" & x(32*32*m*8+865*8+7 downto 32*32*m*8+864*8) & "00000000" & x(32*32*m*8+833*8+7 downto 32*32*m*8+832*8) & "00000000";
                when "1110000000" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= x(32*32*m*8+929*8+7 downto 32*32*m*8+928*8) & "00000000" & x(32*32*m*8+897*8+7 downto 32*32*m*8+896*8) & "00000000" & x(32*32*m*8+865*8+7 downto 32*32*m*8+864*8) & "00000000";
                when "1110100000" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= x(32*32*m*8+961*8+7 downto 32*32*m*8+960*8) & "00000000" & x(32*32*m*8+929*8+7 downto 32*32*m*8+928*8) & "00000000" & x(32*32*m*8+897*8+7 downto 32*32*m*8+896*8) & "00000000";
                when "1111000000" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= x(32*32*m*8+993*8+7 downto 32*32*m*8+992*8) & "00000000" & x(32*32*m*8+961*8+7 downto 32*32*m*8+960*8) & "00000000" & x(32*32*m*8+929*8+7 downto 32*32*m*8+928*8) & "00000000";

                when "0000111111" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= "00000000" & x(32*32*m*8+95*8+7 downto 32*32*m*8+94*8) & "00000000" & x(32*32*m*8+63*8+7 downto 32*32*m*8+62*8) & "00000000" & x(32*32*m*8+31*8+7 downto 32*32*m*8+30*8);--p5 the right edge
                when "0001011111" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= "00000000" & x(32*32*m*8+127*8+7 downto 32*32*m*8+126*8) & "00000000" & x(32*32*m*8+95*8+7 downto 32*32*m*8+94*8) & "00000000" & x(32*32*m*8+63*8+7 downto 32*32*m*8+62*8);
                when "0001111111" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= "00000000" & x(32*32*m*8+159*8+7 downto 32*32*m*8+158*8) & "00000000" & x(32*32*m*8+127*8+7 downto 32*32*m*8+126*8) & "00000000" & x(32*32*m*8+95*8+7 downto 32*32*m*8+94*8);
                when "0010011111" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= "00000000" & x(32*32*m*8+191*8+7 downto 32*32*m*8+190*8) & "00000000" & x(32*32*m*8+159*8+7 downto 32*32*m*8+158*8) & "00000000" & x(32*32*m*8+127*8+7 downto 32*32*m*8+126*8);
                when "0010111111" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= "00000000" & x(32*32*m*8+223*8+7 downto 32*32*m*8+222*8) & "00000000" & x(32*32*m*8+191*8+7 downto 32*32*m*8+190*8) & "00000000" & x(32*32*m*8+159*8+7 downto 32*32*m*8+158*8);
                when "0011011111" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= "00000000" & x(32*32*m*8+255*8+7 downto 32*32*m*8+254*8) & "00000000" & x(32*32*m*8+223*8+7 downto 32*32*m*8+222*8) & "00000000" & x(32*32*m*8+191*8+7 downto 32*32*m*8+190*8);
                when "0011111111" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= "00000000" & x(32*32*m*8+287*8+7 downto 32*32*m*8+286*8) & "00000000" & x(32*32*m*8+255*8+7 downto 32*32*m*8+254*8) & "00000000" & x(32*32*m*8+223*8+7 downto 32*32*m*8+222*8);
                when "0100011111" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= "00000000" & x(32*32*m*8+319*8+7 downto 32*32*m*8+318*8) & "00000000" & x(32*32*m*8+287*8+7 downto 32*32*m*8+286*8) & "00000000" & x(32*32*m*8+255*8+7 downto 32*32*m*8+254*8);
                when "0100111111" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= "00000000" & x(32*32*m*8+351*8+7 downto 32*32*m*8+350*8) & "00000000" & x(32*32*m*8+319*8+7 downto 32*32*m*8+318*8) & "00000000" & x(32*32*m*8+287*8+7 downto 32*32*m*8+286*8);
                when "0101011111" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= "00000000" & x(32*32*m*8+383*8+7 downto 32*32*m*8+382*8) & "00000000" & x(32*32*m*8+351*8+7 downto 32*32*m*8+350*8) & "00000000" & x(32*32*m*8+319*8+7 downto 32*32*m*8+318*8);
                when "0101111111" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= "00000000" & x(32*32*m*8+415*8+7 downto 32*32*m*8+414*8) & "00000000" & x(32*32*m*8+383*8+7 downto 32*32*m*8+382*8) & "00000000" & x(32*32*m*8+351*8+7 downto 32*32*m*8+350*8);
                when "0110011111" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= "00000000" & x(32*32*m*8+447*8+7 downto 32*32*m*8+446*8) & "00000000" & x(32*32*m*8+415*8+7 downto 32*32*m*8+414*8) & "00000000" & x(32*32*m*8+383*8+7 downto 32*32*m*8+382*8);
                when "0110111111" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= "00000000" & x(32*32*m*8+479*8+7 downto 32*32*m*8+478*8) & "00000000" & x(32*32*m*8+447*8+7 downto 32*32*m*8+446*8) & "00000000" & x(32*32*m*8+415*8+7 downto 32*32*m*8+414*8);
                when "0111011111" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= "00000000" & x(32*32*m*8+511*8+7 downto 32*32*m*8+510*8) & "00000000" & x(32*32*m*8+479*8+7 downto 32*32*m*8+478*8) & "00000000" & x(32*32*m*8+447*8+7 downto 32*32*m*8+446*8);
                when "0111111111" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= "00000000" & x(32*32*m*8+543*8+7 downto 32*32*m*8+542*8) & "00000000" & x(32*32*m*8+511*8+7 downto 32*32*m*8+510*8) & "00000000" & x(32*32*m*8+479*8+7 downto 32*32*m*8+478*8);
                when "1000011111" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= "00000000" & x(32*32*m*8+575*8+7 downto 32*32*m*8+574*8) & "00000000" & x(32*32*m*8+543*8+7 downto 32*32*m*8+542*8) & "00000000" & x(32*32*m*8+511*8+7 downto 32*32*m*8+510*8);
                when "1000111111" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= "00000000" & x(32*32*m*8+607*8+7 downto 32*32*m*8+606*8) & "00000000" & x(32*32*m*8+575*8+7 downto 32*32*m*8+574*8) & "00000000" & x(32*32*m*8+543*8+7 downto 32*32*m*8+542*8);
                when "1001011111" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= "00000000" & x(32*32*m*8+639*8+7 downto 32*32*m*8+638*8) & "00000000" & x(32*32*m*8+607*8+7 downto 32*32*m*8+606*8) & "00000000" & x(32*32*m*8+575*8+7 downto 32*32*m*8+574*8);
                when "1001111111" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= "00000000" & x(32*32*m*8+671*8+7 downto 32*32*m*8+670*8) & "00000000" & x(32*32*m*8+639*8+7 downto 32*32*m*8+638*8) & "00000000" & x(32*32*m*8+607*8+7 downto 32*32*m*8+606*8);
                when "1010011111" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= "00000000" & x(32*32*m*8+703*8+7 downto 32*32*m*8+702*8) & "00000000" & x(32*32*m*8+671*8+7 downto 32*32*m*8+670*8) & "00000000" & x(32*32*m*8+639*8+7 downto 32*32*m*8+638*8);
                when "1010111111" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= "00000000" & x(32*32*m*8+735*8+7 downto 32*32*m*8+734*8) & "00000000" & x(32*32*m*8+703*8+7 downto 32*32*m*8+702*8) & "00000000" & x(32*32*m*8+671*8+7 downto 32*32*m*8+670*8);
                when "1011011111" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= "00000000" & x(32*32*m*8+767*8+7 downto 32*32*m*8+766*8) & "00000000" & x(32*32*m*8+735*8+7 downto 32*32*m*8+734*8) & "00000000" & x(32*32*m*8+703*8+7 downto 32*32*m*8+702*8);
                when "1011111111" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= "00000000" & x(32*32*m*8+799*8+7 downto 32*32*m*8+798*8) & "00000000" & x(32*32*m*8+767*8+7 downto 32*32*m*8+766*8) & "00000000" & x(32*32*m*8+735*8+7 downto 32*32*m*8+734*8);
                when "1100011111" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= "00000000" & x(32*32*m*8+831*8+7 downto 32*32*m*8+830*8) & "00000000" & x(32*32*m*8+799*8+7 downto 32*32*m*8+798*8) & "00000000" & x(32*32*m*8+767*8+7 downto 32*32*m*8+766*8);
                when "1100111111" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= "00000000" & x(32*32*m*8+863*8+7 downto 32*32*m*8+862*8) & "00000000" & x(32*32*m*8+831*8+7 downto 32*32*m*8+830*8) & "00000000" & x(32*32*m*8+799*8+7 downto 32*32*m*8+798*8);
                when "1101011111" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= "00000000" & x(32*32*m*8+895*8+7 downto 32*32*m*8+894*8) & "00000000" & x(32*32*m*8+863*8+7 downto 32*32*m*8+862*8) & "00000000" & x(32*32*m*8+831*8+7 downto 32*32*m*8+830*8);
                when "1101111111" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= "00000000" & x(32*32*m*8+927*8+7 downto 32*32*m*8+926*8) & "00000000" & x(32*32*m*8+895*8+7 downto 32*32*m*8+894*8) & "00000000" & x(32*32*m*8+863*8+7 downto 32*32*m*8+862*8);
                when "1110011111" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= "00000000" & x(32*32*m*8+959*8+7 downto 32*32*m*8+958*8) & "00000000" & x(32*32*m*8+927*8+7 downto 32*32*m*8+926*8) & "00000000" & x(32*32*m*8+895*8+7 downto 32*32*m*8+894*8);
                when "1110111111" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= "00000000" & x(32*32*m*8+991*8+7 downto 32*32*m*8+990*8) & "00000000" & x(32*32*m*8+959*8+7 downto 32*32*m*8+958*8) & "00000000" & x(32*32*m*8+927*8+7 downto 32*32*m*8+926*8);
                when "1111011111" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= "00000000" & x(32*32*m*8+1023*8+7 downto 32*32*m*8+1022*8) & "00000000" & x(32*32*m*8+991*8+7 downto 32*32*m*8+990*8) & "00000000" & x(32*32*m*8+959*8+7 downto 32*32*m*8+958*8);

                when "1111100000" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= "000000000000000000000000" & x(32*32*m*8+993*8+7 downto 32*32*m*8+992*8) & "00000000" & x(32*32*m*8+961*8+7 downto 32*32*m*8+960*8) & "00000000";--p6 the left bottom corner

                when "1111100001" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= "000000000000000000000000" & x(32*32*m*8+994*8+7 downto 32*32*m*8+992*8) & x(32*32*m*8+962*8+7 downto 32*32*m*8+960*8);--p7 the bottom edge
                when "1111100010" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= "000000000000000000000000" & x(32*32*m*8+995*8+7 downto 32*32*m*8+993*8) & x(32*32*m*8+963*8+7 downto 32*32*m*8+961*8);
                when "1111100011" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= "000000000000000000000000" & x(32*32*m*8+996*8+7 downto 32*32*m*8+994*8) & x(32*32*m*8+964*8+7 downto 32*32*m*8+962*8);
                when "1111100100" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= "000000000000000000000000" & x(32*32*m*8+997*8+7 downto 32*32*m*8+995*8) & x(32*32*m*8+965*8+7 downto 32*32*m*8+963*8);
                when "1111100101" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= "000000000000000000000000" & x(32*32*m*8+998*8+7 downto 32*32*m*8+996*8) & x(32*32*m*8+966*8+7 downto 32*32*m*8+964*8);
                when "1111100110" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= "000000000000000000000000" & x(32*32*m*8+999*8+7 downto 32*32*m*8+997*8) & x(32*32*m*8+967*8+7 downto 32*32*m*8+965*8);
                when "1111100111" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= "000000000000000000000000" & x(32*32*m*8+1000*8+7 downto 32*32*m*8+998*8) & x(32*32*m*8+968*8+7 downto 32*32*m*8+966*8);
                when "1111101000" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= "000000000000000000000000" & x(32*32*m*8+1001*8+7 downto 32*32*m*8+999*8) & x(32*32*m*8+969*8+7 downto 32*32*m*8+967*8);
                when "1111101001" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= "000000000000000000000000" & x(32*32*m*8+1002*8+7 downto 32*32*m*8+1000*8) & x(32*32*m*8+970*8+7 downto 32*32*m*8+968*8);
                when "1111101010" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= "000000000000000000000000" & x(32*32*m*8+1003*8+7 downto 32*32*m*8+1001*8) & x(32*32*m*8+971*8+7 downto 32*32*m*8+969*8);
                when "1111101011" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= "000000000000000000000000" & x(32*32*m*8+1004*8+7 downto 32*32*m*8+1002*8) & x(32*32*m*8+972*8+7 downto 32*32*m*8+970*8);
                when "1111101100" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= "000000000000000000000000" & x(32*32*m*8+1005*8+7 downto 32*32*m*8+1003*8) & x(32*32*m*8+973*8+7 downto 32*32*m*8+971*8);
                when "1111101101" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= "000000000000000000000000" & x(32*32*m*8+1006*8+7 downto 32*32*m*8+1004*8) & x(32*32*m*8+974*8+7 downto 32*32*m*8+972*8);
                when "1111101110" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= "000000000000000000000000" & x(32*32*m*8+1007*8+7 downto 32*32*m*8+1005*8) & x(32*32*m*8+975*8+7 downto 32*32*m*8+973*8);
                when "1111101111" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= "000000000000000000000000" & x(32*32*m*8+1008*8+7 downto 32*32*m*8+1006*8) & x(32*32*m*8+976*8+7 downto 32*32*m*8+974*8);
                when "1111110000" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= "000000000000000000000000" & x(32*32*m*8+1009*8+7 downto 32*32*m*8+1007*8) & x(32*32*m*8+977*8+7 downto 32*32*m*8+975*8);
                when "1111110001" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= "000000000000000000000000" & x(32*32*m*8+1010*8+7 downto 32*32*m*8+1008*8) & x(32*32*m*8+978*8+7 downto 32*32*m*8+976*8);
                when "1111110010" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= "000000000000000000000000" & x(32*32*m*8+1011*8+7 downto 32*32*m*8+1009*8) & x(32*32*m*8+979*8+7 downto 32*32*m*8+977*8);
                when "1111110011" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= "000000000000000000000000" & x(32*32*m*8+1012*8+7 downto 32*32*m*8+1010*8) & x(32*32*m*8+980*8+7 downto 32*32*m*8+978*8);
                when "1111110100" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= "000000000000000000000000" & x(32*32*m*8+1013*8+7 downto 32*32*m*8+1011*8) & x(32*32*m*8+981*8+7 downto 32*32*m*8+979*8);
                when "1111110101" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= "000000000000000000000000" & x(32*32*m*8+1014*8+7 downto 32*32*m*8+1012*8) & x(32*32*m*8+982*8+7 downto 32*32*m*8+980*8);
                when "1111110110" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= "000000000000000000000000" & x(32*32*m*8+1015*8+7 downto 32*32*m*8+1013*8) & x(32*32*m*8+983*8+7 downto 32*32*m*8+981*8);
                when "1111110111" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= "000000000000000000000000" & x(32*32*m*8+1016*8+7 downto 32*32*m*8+1014*8) & x(32*32*m*8+984*8+7 downto 32*32*m*8+982*8);
                when "1111111000" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= "000000000000000000000000" & x(32*32*m*8+1017*8+7 downto 32*32*m*8+1015*8) & x(32*32*m*8+985*8+7 downto 32*32*m*8+983*8);
                when "1111111001" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= "000000000000000000000000" & x(32*32*m*8+1018*8+7 downto 32*32*m*8+1016*8) & x(32*32*m*8+986*8+7 downto 32*32*m*8+984*8);
                when "1111111010" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= "000000000000000000000000" & x(32*32*m*8+1019*8+7 downto 32*32*m*8+1017*8) & x(32*32*m*8+987*8+7 downto 32*32*m*8+985*8);
                when "1111111011" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= "000000000000000000000000" & x(32*32*m*8+1020*8+7 downto 32*32*m*8+1018*8) & x(32*32*m*8+988*8+7 downto 32*32*m*8+986*8);
                when "1111111100" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= "000000000000000000000000" & x(32*32*m*8+1021*8+7 downto 32*32*m*8+1019*8) & x(32*32*m*8+989*8+7 downto 32*32*m*8+987*8);
                when "1111111101" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= "000000000000000000000000" & x(32*32*m*8+1022*8+7 downto 32*32*m*8+1020*8) & x(32*32*m*8+990*8+7 downto 32*32*m*8+988*8);
                when "1111111110" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= "000000000000000000000000" & x(32*32*m*8+1023*8+7 downto 32*32*m*8+1021*8) & x(32*32*m*8+991*8+7 downto 32*32*m*8+989*8);

                when "1111111111" => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= "00000000000000000000000000000000" & x(32*32*m*8+1023*8+7 downto 32*32*m*8+1022*8) & "00000000" & x(32*32*m*8+991*8+7 downto 32*32*m*8+990*8);--p8 the right bottom corner

                when others => x_single(3*3*m*8+3*3*8-1 downto 3*3*m*8) <= x((32*32*m+I+33)*8+7 downto (32*32*m+I+31)*8) & x((32*32*m+I+1)*8+7 downto (32*32*m+I-1)*8) & x((32*32*m+I-31)*8+7 downto (32*32*m+I-33)*8);--p4 the center part
            end case;
        end process;
    end generate;

    process(S, x)
    begin
        case to_integer(unsigned(S)) is
            when 0 => c <= "0000";--p0
            when 1 to 30 => c <= "0100";--p1
            when 31 => c <= "0001";--p2
            when 32 | 64 | 96 | 128 | 160 | 192 | 224 | 256 | 288 | 320 | 352 | 384 | 416 | 448 | 480 | 512 | 544 | 576 | 608 | 640 | 672 | 704 | 736 | 768 | 800 | 832 | 864 | 896 | 928 | 960 => c <= "0101"; --p3
            when 63 | 95 | 127 | 159 | 191 | 223 | 255 | 287 | 319 | 351 | 383 | 415 | 447 | 479 | 511 | 543 | 575 | 607 | 639 | 671 | 703 | 735 | 767 | 799 | 831 | 863 | 895 | 927 | 959 | 991 => c <= "0110"; --p5
            when 992 => c <= "0010"; --p6
            when 993 to 1022 => c <= "0111"; --p7
            when 1023 => c <= "0011"; --p8
            when others => c <= "1000"; --p4
        end case;
    end process;
end Behavioral;
