library IEEE;
use IEEE.Std_logic_1164.all;
use IEEE.Numeric_Std.all;
use IEEE.STD_LOGIC_TEXTIO.ALL;
library STD;
use STD.TEXTIO.ALL;
use std.env.all; -- VHDL 2008

entity single_step_fc_tb is
end;

architecture bench of single_step_fc_tb is

  component single_step_fc
      generic (
          x_width: integer;
          z_width: integer
      );
      port (
          x : in STD_LOGIC_VECTOR(x_width-1 downto 0);
          w : in STD_LOGIC_VECTOR(x_width-1 downto 0);
          z : out STD_LOGIC_VECTOR(z_width-1 downto 0)
      );
  end component;

  signal x: STD_LOGIC_VECTOR(8192-1 downto 0);
  signal w: STD_LOGIC_VECTOR(8192-1 downto 0);
  signal z: STD_LOGIC_VECTOR(14 downto 0) ;

begin

  -- Insert values for generic parameters !!
  uut: single_step_fc generic map ( x_width => 8192,
                                    z_width =>15  )
                         port map ( x       => x,
                                    w       => w,
                                    z       => z );

  stimulus: process
  begin
  
    -- Put initialisation code here
    w <= "11101101011110001100110101111111100110111001011001111011100010001010000010001001110001011100000001100011001111111111111110000011011001111111000110111001001110111011110000000100111011100110101011000100011101110110111101110001001101110100110000000101111110111011111100111011110100000111000000100010110110110110111111011111101101010110100011110001110111110100111101010010110101111011111100000001000011101010001110101111111100001010100110000100010111101001100111111011101101100010010011101000000111111111111111101110100000000100000000100001011010100100111111111011101000001010111011110110111101110100110001101110110011110111111111010101001101011111011010110001010100110010000001111111111111111111010111100111010100000010000010110110000011011111110111111101010001001100111001110111101111011011000000000111111101100111000010000101111111111001011001101111001100110011000110010111001111111011011000111111110111011000110100011101001001110100011111001000001101010000001111000111110010010100101000100101011111111110001000101111101110011111000010100111010001001101100011110000000100000101010100000011001101110011011101100000001100000111010011010001001011101111100111011011100110010101011111011101011101100000000101100110111000011001100000101001011000010011110101111000010111111111111001100111100101001111111011101001010101100011111001111111000110010000111001001011110111111100111110010011000010011000100010011001111001011000000111100101110101101100110101111111110111100011111110111111010011111111101101000000110100010100000100000000000100001001010101001110101010111111110111111111101011110010111100100000000000110100010000001010011100000100111011000010011001101100000000101000001001101110100001111100111001101101000000001011111001100101100111000111111111111101000011110101110101000110101111100101100110011101111001110110110101101101101110101111111111111100110101011111101000001000100111101011000001111010100001101111110011110110000110100111010111110010000001100011011111111101110101100101110101110011110000010011010011010110110110001101111100001110000000000111011000000000100011100010011001111101011111001011011010000100000000101000100100111101010101101111111110111000000010101101101011101111000001111101100110001000011011011110000011011110111001011110001111011111111000001100011011100000011001111111111011000010111010001111000011010111000100001110100101110111000111111001000110111001111010111100001101111001110101100110000110101110000011110111001111111111110000110100100000001101011111111111101001001000010010100111110111010011100101000000100110000101101110100000011100001001101100110101011111101110101011100000111111001111110000010000110011101001101111101010001010010110100100000001010000110001100001000011011000110100001000011110010000000001100001000100000001100101111100000101110010010001010101010001101110110111100101100100110110111010001011111101111110101111100010000000010000101000101110001010101000101111110010000111101110000100111001000000101100010110001110001000111110111111011011100000010101010001100001111101100110000010000001001111111011111100111000001100011100111110110010110011111100001101011011101111000010111001010101101111101111100010110001100000100111000000010100010111000011110001111000011110000110101101100110011010010011101111100001101111100110110000000100111000010100011001110101110010100110001101011110110110001111010101011111101111101101010000011011100000001011110101001101010001100011110111001011001010000010011100000001101011101001111010011000010001001111111001101100010101101110110010011110110110001101110110100100101110011111000011011100001010000000011111010000110000010100100010000101110101001011111110000010101111111101111001011101100010011011001101100011110111100010010011101111000101100111010100011110111101111110111111001101011100100100000110111101111111111111001110111111101011101110100011111000110101011111110110001100111010000000010111110101010010001111111111111000100111000100110010110101100110111110111110011100100011000000001001010101010100110100000110101111100101110011111010111101001111100100101110000111011010100111110110111000001010111010011001001010110011101000101011110000001011010101101000000111000001000000111111011111110010100111010110111011111010111101111101111111000100110011101011100001100110111011010011001011100001111101101111101111110000100000001110101001101111011110101111000110110110000100101100101100001110111101100001001010111101001000010110111110101111110111111011100100100101100111000001011111011001000100000011111100101111111001000001010001111110101101010001111110000100110010011011010101000000000111000111011101101010000011110111111100101001010100001011000001011110011110100100011011100010111101111111111001101101011111000011010111111101011110011111011111111001101111000001100110001100100101011000001011111001000001100111101111101100111110010110100010110011101101000011001111000001101100111111111110111010111110110101100011110000100111101110101110001001000001100010101010111010101110001110101011010001101011111000011111111001111110111011011011000100111111111101001000000000010000001100111111011011110001011111110011101001111100000000111111111101010100111101111110000001110111100111111100100000000000001001000111000010110010000100000000101111010001111100101110001111011011100001100110100011100100100011110011011000111000110101111111001111011100010010101010101101111110001101100001101001101111110110011101101101011100000001101110110111011011101011011101101100110111010001111111001101110011100011011100111111001011001010010101111011100110111111100111010001101011011111111010000001100101110100000101110111111010001001100110001010110000001001110101111110101101010101011011111111111111010101011001010111100010100010001000011101001100010100010010110000101101000011100011001000010111101100100101101111111000010110111000100000011011001001011001000000010100101101010111001000111010000111111011110000010101001001110111011110101010010101001011111001111110110110111110011100011000000100101011100000111000010110000000110000111011001101001110000100110100101101101110110011111111111010111011111111001110011011010011111110110100011100110101111111110000000001001011101011110111111100101001011111111111000011101101110001011100010100010101001001000111000011100001001011100010110100100000111011010110001111100000011100000110011111111000100000011011000111000000111001111111110010101111110110000110101111110111011111111101011111101011110111100100111111111101110011010110101010011111100100001001010100001010011101100111100110111011011111010001100001000101101001100000111010011001001001110001111011100010101101001110110011010100000001110101000001000000000110101100011010000110000111111001111011000111010101101000101111001110101011100011111001111011111100011111111011011100010111101110100001100100110011000100110111100110011110011110110001010101111011001001011111100011010000011111011111011010001010001000110011110000111101111110011100011100111111011001110010101101100101100111111111001010001011111101100001000001110101011110101010000101100111110000100010010001110011111110101001111100100011010011000111000011010011001110010110110010010101110101100010011100011100101101100011110110100100001101001011111001010111111100100001001001110111011111001100110101111100011000110101001100011010010011011001010111000000101101111110000001111000110001000110100100100011111010100000100111101001011010111110100011100001101001101100010010111001100101111110101101000010000010111000111110110011100110001111100111001001100000000111111101110111110110001000101111011110100010100110010001011111101101101001011100101110110001011001111000011100001110110010010000011000001111000011011111010110001010000010001000111111000101011111000111010110111101100000011111110110011101101101110010011101011111001110010111011100110000011110010101001000111011011101111111010000010101001110101101000110100101100111000111101010010100010000101001011000011100100101000010001011100110010111011010001100100100001000010000110010110010010111111010001010110100001001101101111001100101101111111111011111001111111010011111111110110000000111000011000010011101111100010101101111110001010110110011100101111010101000110000100110110011111011110001101010101101111100010000111110101101000010011110010001000110010111000001111000";
    x <= "00101110111011110110010001000001111111010001001010111101101100010000000000000000000000000000000001100000000010000100001000100000000000100000010011100101010010101100010000101011111111111111111000000001000011000000011000100000000101010110000100100101111010111111111111111111000000000100010001110111111111110010010000000000111111111111111100000100011100010000000000000000111111011111111111110111000100011111010011110011000000010000000000000000010000000010001000100100100000100110100011111111111111111100110011110011000000100100000000000000001000001100111001111000000000001000000010000010001000000000001101010100111111110111111110011011001000110000000000001100000100000010100000010000010101000101010011100001000000000000010000000010010000001011111111111111000100010101010011001010001010001110000011001011100000100000000000000001010100001111111111111011000000000011000010000100000100000100001000000000011000000000000000000011110001110000000101010000000000001000001011111111111111111000001000000000000001110101000000000000001101001011000100111110000000000000000000010000010100010000000000000000010001001000000010111111111111111000010001000001000000000000000000100010000001000000001000000110010001000000000000000010111001011111001101001100111111111111111111110111111111010010001000101000010000000110010000100010010011000000001001000000011111000011000011110001111111100000000000000000000001001000000000111111111011100000000000000000000000000000000011110000001010000000111001100001101000100101010011111111111111110011100100100000111111111111111100100000110000010000000100100000111001001001100100000010000000001101010100011111111111111011101111111111111111110111001011101111000000000100000001000100011100000000000000001010100001010100001000000100010010011111111111111111011111111111111100000000000000001000011000101011111111111111111100000000010010000001000100000000100000100010011000000000100000111111111111111111001000000000010011111111111111110000011001000000100001101100000000000000000000001100100000110010000000000100000011000100101101001111101110101111100001010100000101111111111111110000010011000000111101111111111100011010001010010000010011101100000000000000000000000000000000001111000011110111010010000110000001000111000101000010111111001010100011111101100111111111011111110000011001000000111111111111111001111111001011000011000000000000000001000111001011111111110111011001001111111111000000000100000111111111001111111111111111111111000000000000000001001110111000010000100000000000000000100000000010000000000000000000001000000000010111111111101111110001000111110100010100000000111111111111111100000000000000000000000000000000001000110101111100000000000000000100010000000000000000000100000011111001000111110110000100100001000001000000010011111011000011100000000000000000010000001100000111111111111111110001000000000000011100100000000111111111111111110000000000000001000001000010000000100010011010111100100010010001001000000101011000000101000010011000011100000000001000100000000000000000101000001011111111111111111111111011101111111111111111110000000000000000111111111111111100000000000000000000101000000000001111011001101100100001000000000000010000000000000000000000000000000011000000101101101101111110111000001001000001100100001000010000011000000010000000000000001000000010001101001111111111111111010010100011001110110101111001111111111111111111001000000000000111111111101111110010001001000000000000100110001000110011001111011011011011111101111011111101111100010010100001001101110110011111000000100000000011110111111111010000000100000000000110100000000011101100100000000000001000000000000011001100101101000000000010001111111111111111110110111111111101110111111111111111111011010111111110111111111100100001000001001111111111111111000000000000000110111111101111010010000010110000101101111011111100001101111110001011111111111111100000100000100010000010010000000010000100010000000000000010000000000000001000000011001011101111111111111111111110111000001000011100000000010110000000000000000000000001000010100011100101011110100000100000000001111111111110110000010101000000011100000001000000000001001100000111011000000110100010100000000001000010000100000011111101011111000000100000000010111011111111011101100100001111010000000000000011111111111111110000001011101100000111111111111100001110100110011111111111111111000001010101101111011111001110111111111100111110000001101100100111111101111111110111001010001010001000100010000000000000000000001111110111111111000001010101100011111101001111110000000011100010111111101111111101000000001100000000000000000001000000100001000001011100101100010000001000000000010011101101010010000010000000001111001111111111010000001011000100000000010100000010011011111011111111111111111111011100111100010111011101111101001000000100011111111011000011110000000000000000110010000010000000110001000000010001101100000000000000001100101000010101000000001000001010100001000000000000000000010010000000001111111110111111001001101110000011110000000110000000010000000000001101111011101011111111111111110000000000101000011101110011000011111111011011111100110111010111001000010010000011111101111111110000000001010000100000000100000001000100000000001111111111111111000000100000000011111011101111111100010100000110100000110000000001110101110000010000001000000000111100110000000000001010100000000000100001000000000000011010000000010100100010000000000010000000111111011111110100100011111011110000100011000000000000000110000001101100101100000000000000000000000000100011000110000010001000000001000000100001000000001010000000010000100000001101010111011111000000010010000000110011111111110011010101100100000000000000000000000000010000001101001110000100011000000001000001001100101101110010000000000000010111000001000011111111111111111101100111101111000001000100000101000000010000001111111110001000001100110011111000000000100000001011110111111111111111111111111111111111111111110000000100000010011101011101101001110000010000010000100010100000000000000000000001100110111011111000001000100000001000000010000000000010010000011111111101111111000000000000000100000000101000000000010011001001000000100110000000000000000000000000110010100101011011000111000100000010101000100001101101111010000000101110100111001011111111111111111110111111111111110101000101001000100100000000000000000000001100000001001000100110000000001111111110011001111100110011011100000110010000010000000010100110111111111111011100010001000000000000010011000000100000010000000000000110001000001111001001010000111110101111110101010001000000010000001000101000111111111111111111111011010110010010011001100000000101000110000101000001001101011100111101011110011111111111101110000010000000011010000001100100000000000000000010000000110001011111111111111111111111111111111100001100100000001100010000010010010000000110000010110111001100010011101011100111000000000100000011111111111111110000001011100000000000100110000010010011111111110000011000000000111111111111111111010010001111001111001110111110000001000000000000000010000010000000011011101101111111111111111100000000000000000000001000000000011000101100001110111111111111110001101011111111000001010010000000000100101000000000001000001000111101111111111100000000000100000000000000110000000001000000000000000010000000000111000011100101000000100010000100000000000000001111111111111111111111111111111111001000100001001111111110011011111111111111111111011001110110110000000000000000000000000000000000000000000000001100100110111100100011110101000100100000000000000011001000100000100000001001000010010010001000110000011100110100011001001110111111110010011111110000000000000000010101110011000000000000000000001111111111011111111111111111111100000000000000010000000000000110000000000000100100000010000000101000001100000000011101101101101110000101010100000110000000100100111111111111111100000000001000000000001011000100000000000100100001000110001000001000010011011111001100010010000000000000000000000011001011100000000110001011110000100000010000000000001000000001000000000010000000000000011000001111111011110111010000101000000011111111111111110000011000000000010000000000001011111110111111111111100001000110111001111011111100110110110010001100010110001111000000000000000000100010001000000000000000100000";
    
    

    -- Put test bench stimulus code here

    wait;
  end process;
  process(z)
    variable tmp_int : integer; --STD_LOGIC_VECTOR(4*4*512-1 downto 0);
    variable tmp_line : line;
    
  begin
    tmp_int := to_integer(signed(z));
    write(tmp_line, tmp_int);
    writeline(output, tmp_line);
  end process;


end;